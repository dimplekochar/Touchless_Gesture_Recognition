receiver ir
.include ua741.txt
Is 1 2 dc 200u
vdc 1 0 dc 5
r1 2 3 10k
X1 0 3 5 6 7 ua741
vdd 5 0 dc 15
vss 6 0 dc -15
r2 5 7 100k
r3 7 8 1k
X2 0 8 5 6 11 ua741
r4 8 11 10k
.tran 0.0001 10ms
.control
run
plot v(11)
.endc
.end
 


receiver
.include Diode_1N914.txt
.include lm324.txt
X1 11 12 1 0 13 LM324
X2 11 22 1 0 23 LM324
X3 11 32 1 0 33 LM324
X4 33 42 1 0 42 LM324
X5 51 11 1 0 53 LM324
vss 1 0 dc 12
r1 2 3 10k
c1 3 12 10n
r2 1 11 1k
r3 11 0 1k
c2 11 0 1u
c3 11 0 0.22u
r4 12 13 62k
r5 13 4 2.2k
r6 4 11 1k
c4 4 22 1n
c5 4 23 1n
r7 22 23 15.45k
c6 22 23 12p
r8 23 5 10k
c7 5 32 10n
r9 32 33 75k
d1 42 51 1N914
r10 51 0 61.6k
c8 51 0 2n
r11 53 6 12k
r12 6 0 10k
vin 2 0 sin(0 9m 40k) 
.tran 0.0001 0.5ms
.control
run
plot v(6)
.endc
.end

